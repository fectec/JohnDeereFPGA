LIBRARY	IEEE;
USE	IEEE.STD_LOGIC_1164.ALL;

ENTITY Decoder_BCDTo7Seg IS

	PORT	(	
				BCD		:	IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
				Segments	:	OUT	STD_LOGIC_VECTOR(13 DOWNTO 0)
		);
			
END ENTITY Decoder_BCDTo7Seg;

ARCHITECTURE Dataflow of Decoder_BCDTo7Seg IS 
		
BEGIN

	Segments 	<= 	"10000001000000" 	WHEN 	BCD = "0000" 	ELSE	-- 0
				"10000001111001" 	WHEN 	BCD = "0001" 	ELSE	-- 1
				"10000000100100" 	WHEN 	BCD = "0010" 	ELSE	-- 2
				"10000000110000" 	WHEN 	BCD = "0011" 	ELSE	-- 3
				"10000000011001" 	WHEN 	BCD = "0100" 	ELSE	-- 4
				"10000000010010" 	WHEN 	BCD = "0101" 	ELSE	-- 5
				"10000000000010" 	WHEN 	BCD = "0110" 	ELSE	-- 6
				"10000001111000" 	WHEN 	BCD = "0111" 	ELSE	-- 7
				"10000000000000" 	WHEN 	BCD = "1000" 	ELSE	-- 8
				"10000000010000" 	WHEN 	BCD = "1001" 	ELSE	-- 9
				"11110011000000" 	WHEN 	BCD = "1010" 	ELSE	-- 10 
				"11110011111001" 	WHEN 	BCD = "1011" 	ELSE	-- 11
				"11110010100100" 	WHEN 	BCD = "1100" 	ELSE	-- 12
				"11110010110000" 	WHEN 	BCD = "1101" 	ELSE	-- 13
				"11110010011001" 	WHEN 	BCD = "1110" 	ELSE	-- 14
				"11110010010010" 	WHEN 	BCD = "1111"; 		-- 15

END ARCHITECTURE Dataflow;
